folded_cascode_amp test

.include "../../../pdk/gf180/ngspice/design.ngspice"

.lib "../../../pdk/gf180/ngspice/sm141064.ngspice" sf


.param wp11=1.0e-6 lp11=300.0e-9 mp11=1
.param wp10=1.0e-6 lp10=300.0e-9 mp10=1
.param  wp7=9.9334e-05 lp7=300.0e-9  mp7=1
.param  wp6=4.9157e-05 lp6=300.0e-9  mp6=1
.param  wp9=1.0e-6 lp9=300.0e-9  mp9=1
.param wn13=5.0e-7 ln13=300.0e-9 mn13=1
.param wn15=1.0e-6 ln15=300.0e-9 mn15=1
.param wn21=9.9165e-05 ln21=300.0e-9 mn21=1
.param c1=10p
.param c2=10p
.param ibias=30u
.param vddh=3.6
.param vcm=0.5*vddh
.param vtran=0.22*vddh

* for transient simulation
.PARAM val0 = 'vtran-0.15'
.PARAM val1 = 'vtran+0.15'
.PARAM GBW_ideal = 5e4
.PARAM STEP_TIME = '10/GBW_ideal'



* Cell name: Folded_cascode
.subckt Folded_cascode gnda vdda vinn vinp vout
xm11 VOUT net050 VDDA VDDA pmos_3p3   l=lp11 w=wp11 m=mp11
xm7 net043 net013 VDDA VDDA pmos_3p3  l=lp7 w=wp7 m=mp7
xm10 net013 net050 VDDA VDDA pmos_3p3 l=lp10 w=wp10 m=mp10
xm6 net050 VOUTN VDDA VDDA pmos_3p3   l=lp6 w=wp6 m=mp6*8
xm5 VOUTN VOUTN VDDA VDDA pmos_3p3    l=lp6 w=wp6 m=mp6*8
xm9 net063 VINP net31 net31 pmos_3p3  l=lp9 w=wp9 m=mp9
xm8 DM_2 VINN net31 net31 pmos_3p3    l=lp9 w=wp9 m=mp9
xm4 net31 net1 VDDA VDDA pmos_3p3     l=lp6 w=wp6 m=2*mp6
xm3 VB3 net1 VDDA VDDA pmos_3p3       l=lp6 w=wp6 m=mp6
xm2 DM_1 net1 VDDA VDDA pmos_3p3      l=lp6 w=wp6 m=mp6
xm1 VB4 net1 VDDA VDDA pmos_3p3       l=lp6 w=wp6 m=mp6
xm0 net1 net1 VDDA VDDA pmos_3p3      l=lp6 w=wp6 m=mp6
xm59 net013 VB4 GNDA GNDA nmos_3p3    l=ln13 w=wn13 m=mn13*8
xm22 VOUT net043 GNDA GNDA nmos_3p3   l=ln21 w=wn21 m=mn21
xm21 net043 net043 GNDA GNDA nmos_3p3 l=ln21 w=wn21 m=mn21
xm19 DM_2 VB4 GNDA GNDA nmos_3p3      l=ln13 w=wn13 m=mn13*8
xm15 VOUTN VB3 DM_2 GNDA nmos_3p3     l=ln15 w=wn15 m=mn15*1
xm20 net063 VB4 GNDA GNDA nmos_3p3    l=ln13 w=wn13 m=mn13*8
xm16 net050 VB3 net063 GNDA nmos_3p3  l=ln15 w=wn15 m=mn15*1
xm17 net54 VB4 GNDA GNDA nmos_3p3     l=ln13 w=wn13 m=mn13*4
xm14 VB3 VB3 GNDA GNDA nmos_3p3       l=ln13 w=wn13 m=mn13
xm12 VB4 VB3 net54 GNDA nmos_3p3      l=ln13 w=wn13 m=mn13*4
xm18 net56 VB4 GNDA GNDA nmos_3p3     l=ln13 w=wn13 m=mn13*4
xm13 DM_1 VB3 net56 GNDA nmos_3p3     l=ln13 w=wn13 m=mn13*4
* Rfix_dm2 DM_2 0 10G
* Rfix_net1 net1 0 10G
I0 net1 GNDA ibias
C1 net050 net013 {c1}
C0 net063 VOUT {c2}
.ends folded_cascode


* Cell name: Folded_cascode_two_stage_TB
V0 in vss dc=0.0 ac=1.0
E1 vin vref in vss -0.5
E0 vip vref in vss 0.5
V1 vdd 0 dc=vddh ac=0
V2 vss 0 dc=0 ac=0
V6 vref vss dc=vcm ac=0
C0 vo vss 10p
X0 vss vdd vin vip vo Folded_cascode


VVISR visr 0 pulse('val0' 'val1' 1u 1p 1p '1*STEP_TIME' 1)
X1 vss vdd vo1 visr vo1 Folded_cascode
CLoad6 vo1 0 500p

* .meas tran t_rise_edge when v(vo1)=1.7 rise=1
* .meas tran t_rise_ param='t_rise_edge - 1u'
* .meas tran t_rise param='t_rise_ * 1e6'
* .meas tran sr_rise param='0.3 / t_rise'
* .meas tran t_fall_edge when v(vo1)=1.7 fall=1
* .meas tran t_fall_ param='t_fall_edge-1u-STEP_TIME'
* .meas tran t_fall param='t_fall_*1e6'
* .meas tran sr_fall param='0.3/t_fall'



.control
set temp=-40
ac dec 10 1 10G
run
set units=degrees
set wr_vecnames
option numdgt=7
wrdata ac.csv v(vo)
op
wrdata dc.csv i(V1)
dc V0 -0.001 0.001 1e-5
wrdata dc_sweep.csv v(vo)

tran 1u 4.01e-4
wrdata tran.csv v(visr) v(vo1)
.endc

.end