
* Instead just load tt corner which is faster
.param mc_mm_switch=0
.param mc_pr_switch=0
.include "../../../pdk/sky130A/libs.tech/ngspice/corners/ss.spice"
*.include "../../../pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice"


.param W_M1=96.02854725718498
.param L_M1=1.5285361856222153
.param W_M2=W_M1 L_M2=L_M1
.param W_M3=74.26867225766182
.param L_M3=0.5013966262340546
.param W_M4=W_M3 L_M4=L_M3
.param W_M5=93.519849807024
.param L_M5=0.5285611003637314
.param W_pass=36.274210065603256
.param L_pass=0.5104859471321106
.param M_pass=110
.param Vb=0.9194943994283675
.param RFB=476.0
.param CFB=0.88p
.param CL=476p
.param vddh=2.0
.param Vref=1.8
.param IL=10m

Vref Vref GND Vref
.save i(vref)
Vb net1 GND Vb
.save i(vb)
IL Vreg net2 dc IL PULSE(10u IL 0 10n 10n 50u 100u 0)
Vdd Vdd GND ac 1 dc vddh
.save i(vdd)
x1 Vdd Vreg Vref net1 GND Vreg ldo
CL Vreg GND {CL}
Rdummy net2 GND 1 m=1
Vref1 Vref1 GND Vref
.save i(vref1)
Vb1 net3 GND Vb
.save i(vb1)
IL1 Vreg1 GND IL
Vdd1 Vdd1 GND vddh
.save i(vdd1)
x2 Vdd1 net4 Vref1 net3 GND Vreg1 ldo
CL1 Vreg1 GND {CL}
Vprobe2 probe net4 dc 0
.save i(vprobe2)
Vprobe1 probe Vreg1 dc 0 ac 1
.save i(vprobe1)
Iprobe1 GND probe dc 0 ac 0
**** begin user architecture code

**** end user architecture code
**.ends


.subckt ldo Vdd Vfb Vref Vb Vss Vreg
x1 Vdd net1 Vfb Vref Vb Vss diff_pair
XM6 Vreg net1 Vdd Vdd sky130_fd_pr__pfet_g5v0d10v5 L=L_pass W=W_pass nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=M_pass m=M_pass
Cfb net2 Vreg {CFB}
Rfb net2 net1 {RFB}
.ends


.subckt diff_pair Vdd vout vinp vinm Vb Vss
XM1 net1 vinp net2 Vss sky130_fd_pr__nfet_g5v0d10v5 L=L_M1 W=W_M1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vout vinm net2 Vss sky130_fd_pr__nfet_g5v0d10v5 L=L_M2 W=W_M2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 vout net1 Vdd Vdd sky130_fd_pr__pfet_g5v0d10v5 L=L_M3 W=W_M3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net1 Vdd Vdd sky130_fd_pr__pfet_g5v0d10v5 L=L_M4 W=W_M4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 Vb Vss Vss sky130_fd_pr__nfet_g5v0d10v5 L=L_M5 W=W_M5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.control
* save all voltage and current
save all
.options savecurrents 
set filetype=ascii
set units=degrees
set temp=125

* high precision simulation
*.OPTIONS maxord=1
.OPTIONS itl1=200
.OPTIONS itl2=200
.OPTIONS itl4=200

* Loop stability
alter IL1 dc=10u
let runs=2
let run=0

alter @Vprobe1[acmag]=1
alter @Iprobe1[acmag]=0

dowhile run<runs
set run=$&run

ac dec 10 1 10G

alter @Vprobe1[acmag]=0
alter @Iprobe1[acmag]=1

let run=run+1
end

let ip11 = ac1.i(Vprobe1)
let ip12 = ac1.i(Vprobe2)
let ip21 = ac2.i(Vprobe1)
let ip22 = ac2.i(Vprobe2)
let vprb1 = ac1.v(probe)
let vprb2 = ac2.v(probe)

*** Middlebrook
let mb = 1/(vprb1+ip22)-1
*** Tian that is preferred
let av = 1/(1/(2*(ip11*vprb2-vprb1*ip21)+vprb1+ip21)-1)

*plot vdb(mb) vp(mb)
*plot vdb(av) vp(av)

wrdata ldo_tb_loop_gain_minload.txt mag(av) vp(av)

* at max load
reset all
alter IL1 dc=10m
let runs=2
let run=0

alter @Vprobe1[acmag]=1
alter @Iprobe1[acmag]=0

dowhile run<runs
set run=$&run

ac dec 10 1 10G

alter @Vprobe1[acmag]=0
alter @Iprobe1[acmag]=1

let run=run+1
end

let ip11 = ac3.i(Vprobe1)
let ip12 = ac3.i(Vprobe2)
let ip21 = ac4.i(Vprobe1)
let ip22 = ac4.i(Vprobe2)
let vprb1 = ac3.v(probe)
let vprb2 = ac4.v(probe)

*** Middlebrook
let mb = 1/(vprb1+ip22)-1
*** Tian that is preferred
let av = 1/(1/(2*(ip11*vprb2-vprb1*ip21)+vprb1+ip21)-1)

*plot vdb(mb) vp(mb)
*plot vdb(av) vp(av)

wrdata ldo_tb_loop_gain_maxload.txt mag(av) vp(av)

* DC sweep
dc Vdd 1 3 0.01
*plot v(Vdd) v(Vreg)
wrdata ldo_tb_dc.txt v(Vreg)

* Transient analysis with load regulation
* do not miss the space between the square bracket and number
* tran 10n 100u
* plot @Rdummy[i]
* plot Vreg
* wrdata ldo_tb_load_reg.txt Vreg
* wrdata ldo_tb_load_reg_current.txt @Rdummy[i] 

* PSRR with max load
ac dec 10 1 10G
*plot vdb(Vreg)
wrdata ldo_tb_psrr_maxload.txt mag(Vreg) vp(Vreg)

* PSRR with min load
alter IL dc=10u
ac dec 10 1 10G
*plot vdb(Vreg)
wrdata ldo_tb_psrr_minload.txt mag(Vreg) vp(Vreg)

.endc


.GLOBAL GND
.end
